`timescale 1ns / 1ps

module ROM (
    input  [31:0] addr,
    output [31:0] data
);
 
    reg [31:0] rom[0:1023];

    initial begin
        
      $readmemh("code.mem",rom);
    
      // GPO test
        // rom[0] = 32'h400007b7; //li      a5,1073741824(0x4000_0000)
        // rom[1] = 32'h0ff00713; //li      a4,255
        // rom[2] = 32'h00e7a023; //sw      a4,0(a5)

        //rom[x] = 32'b_func7 _rs2  _rs1  _f3 _rd   _opcode; //ADD rd  rs1 rs2

        //R-type test
          // rom[0] = 32'b0000000_00001_00010_000_00110_0110011; //ADD x6 x2 x1 -> 6+3 =9
          // rom[1] = 32'b0100000_00001_00010_000_00111_0110011; //SUB x7 x2 x1 -> 6-3 =3
          // rom[2] = 32'b0000000_00001_00011_001_01000_0110011; //SLL x8 x3 x1 -> 9<<3 =1001000 = 72
          // rom[3] = 32'b0000000_00001_00100_101_01001_0110011; //SRL x9 x4 x1 -> -94709717 >> 3 = '0'{-94709717}
          // rom[4] = 32'b0100000_00001_00100_101_01010_0110011; //SRA x10 x4 x1-> -94709717>>3 = '1'{-94709717}
          // rom[5] = 32'b0000000_00001_00100_010_01011_0110011; //SLT x11 x4 x1-> -94709717<3 = 1
          // rom[6] = 32'b0000000_00001_00100_011_01100_0110011; //SLTU x12 x4 x1-> 4,200,257,579 < 3 = 0
          // rom[7] = 32'b0000000_00010_00001_100_01101_0110011; //XOR x13 x1 x2 -> 0011^0110 = 0101 (5)
          // rom[8] = 32'b0000000_00010_00001_110_01110_0110011; //OR  x14 x1 x2 -> 0011 | 0110 = 0111(7)
          // rom[9] = 32'b0000000_00010_00001_111_01111_0110011; //AND x15 x1 x2 -> 0011 & 0110 = 0010 (2)

        // IL-type test
          //rom[x] = 32'b_imm7       _ rs1 _f3 _rd   _opcode; //
            // rom[4] = 32'b000000000010_00001_010_00011_0000011; // LW x3, x1, 2; -> 3+2번째 주소의 값 읽어라. ram[5] = 50
            // rom[0] = 32'b000000000000_00001_000_00011_0000011; // LB x3, x1, 0; -> x1(0)+0번째 주소의 signed Byte값 읽어라. ram[0] = 32'b10101010_01010101_11111111_"11001100"; "zero-extend"
            // rom[1] = 32'b000000000000_00001_001_00100_0000011; // LH x4, x1, 0; -> x1(0)+0번째 주소의 signed half값 읽어라. ram[0] = 32'b10101010_01010101_"11111111_11001100"; "zero-extend"
            // rom[2] = 32'b000000000000_00001_010_00101_0000011; // LW x5, x1, 0; -> x1(0)+0번째 주소의 Byte값 읽어라. ram[0] = 32'b10101010_01010101_11111111_"11001100";
            // rom[3] = 32'b000000000000_00001_100_00110_0000011; // LBU x6, x1, 0; -> x1(0)+0번째 주소의 unsigned Byte값 읽어라. ram[0] = 32'b10101010_01010101_11111111_"11001100";"MSB extend"
            // rom[4] = 32'b000000000000_00001_101_00111_0000011; // LHU x7, x1, 0; -> x1(0)+0번째 주소의 unsigned Byte값 읽어라. ram[0] = 32'b10101010_01010101_11111111_"11001100"; "MSB extend"
        // I-type test
          //rom[x] = 32'b_imm7        _ rs1 _f3 _rd   _opcode; //
            // rom[0] = 32'b0000000_00001_00010_000_00110_0010011; //ADDI x6  x2 1 -> 6+1 =7
            // rom[1] = 32'b0000000_00001_00001_010_00111_0010011; //SLTI x7  x1 1 -> -94709717 < 1 = 1
            // rom[2] = 32'b0000000_00001_00001_011_01000_0010011; //SLTIU x8  x1 1 -> 4,200,257,579 < 1 = 0
            // rom[3] = 32'b0000000_00001_00010_100_01001_0010011; //XORI x9  x2 1 -> 0110 ^ 0001 = 0111 (7)
            // rom[4] = 32'b0000000_00010_00010_110_01010_0010011; //ORI  x10 x2 2 -> 0110 | 0010 = 0110 (6)
            // rom[5] = 32'b0000000_00010_00010_111_01011_0010011; //ANDI x11 x2 2 -> 0110 & 0010 = 0010 (2)

            // rom[0] = 32'b0000000_00001_00010_000_00110_0010011; //ADDI x6  x2 1 -> 6+1 =7
            // rom[1] = 32'b0000000_00001_00010_010_00111_0010011; //SLTI x7  x2 1 -> 6<1 = 0
            // rom[2] = 32'b0000000_00001_00010_011_01000_0010011; //SLTIU x8  x2 1 -> 6 < 1 = 0
            // rom[3] = 32'b0000000_00001_00010_100_01001_0010011; //XORI x9  x2 1 -> 0110 ^ 0001 = 0111 (7)
            // rom[4] = 32'b0000000_00010_00010_110_01010_0010011; //ORI  x10 x2 2 -> 0110 | 0010 = 0110 (6)
            // rom[5] = 32'b0000000_00010_00010_111_01011_0010011; //ANDI x11 x2 2 -> 0110 & 0010 = 0010 (2)
            
        // IStype test
          //rom[x] = 32'b_imm(7)_shift_ rs1 _f3 _rd   _opcode; //
            // rom[6] = 32'b0000000_00001_00010_001_01100_0010011; //SLLI x12 x1 1 -> 6<<1 =0001100 = 12
            // rom[7] = 32'b0000000_00001_00010_101_01101_0010011; //SRLI x13 x1 1 -> 6>>1 = 3
            // rom[8] = 32'b0100000_00001_00101_101_01110_0010011; //SRAI x14 x1 1 -> 6>>1 = 3

        // S_Type test
          //rom[x] = 32'b_imm[11:5]_rs2_ rs1_func3_imm[4:0] _opcode; //
            // rom[0]  = 32'h0ad00093; // addi	x1, x0,173(b10101101)
            // rom[1]  = 32'h00800113; // li		x2, 8
            // rom[2]  = 32'h002091b3; // SLL		x3, x1, x2
            // rom[3]  = 32'h00402023; // sw		x4, 0(x1)
            // rom[4]  = 32'h00100423; // sb    x1, 8(x0)
            // rom[5]  = 32'h001004a3; // sb    x1, 9(x0)
            // rom[6]  = 32'h00100523; // sb    x1, 10(x0)
            // rom[7]  = 32'h001005a3; // sb    x1, 11(x0)
            // rom[8]  = 32'h00301623; // sh   x3, 12(x0)
            // rom[9]  = 32'h003016a3; // sh   x3, 13(x0)
            // rom[10] = 32'h00301723; // sh   x3, 14(x0)
            // rom[11] = 32'h003017a3; // sh   x3, 15(x0)

            // rom[0] = 32'b_0000000_00001_00010_000_00110_0010011; //ADDI x6  x2 1 -> 6+1 =7
            // rom[0] = 32'h0ad00293; // addi	x5, x0,173(b10101101)
            // rom[1] = 32'h00800093; // li		x1, 8
            // rom[2] = 32'h00129333; // SLL		x6, x5, x1
            // rom[2] = 32'h00f0a023; // sw		a5, 0(x1)
            // rom[3] = 32'h00500223; // sb    x5, 4(x0)
            // rom[4] = 32'h005002a3; // sb    x5, 5(x0)
            // rom[5] = 32'h00500323; // sb    x5, 6(x0)
            // rom[6] = 32'h005003a3; // sb    x5, 7(x0)
            // rom[7]  = 32'h00601423; // sh   x6, 8(x0)
            // rom[8]  = 32'h006014a3; // sh   x6, 9(x0)
            // rom[9]  = 32'h00601523; // sh   x6, 10(x0)
            // rom[10] = 32'h006015a3; // sh   x6, 11(x0)

          // B-type test
            //imm[12]_imm[10:5]_rs2[4:0]_rs1[4:0]_func[2:0]_imm[4:1]_imm[11]_opcode[6:0]
            // rom[0] = 32'h00402083; //LW x1 4(x0)  -> x1 = ram[1] = 1
            // rom[1] = 32'h00002103; //LW x2 0(x0)  -> x2 = ram[0] = 32'hffffffff;
            // rom[2] = 32'b0_000000_00010_00001_000_0100_0_1100011; //BEQ x1, x2, 8  -> 1==ffff -> 거짓. (다음에 값나옴)
            // rom[3] = 32'b00000000000000000000_00011_0010111; //AUIPC x3 0 -> RF[3] = PC(0x0c) 
            // rom[4] = 32'b0_000000_00010_00001_001_0100_0_1100011; //BNE x1, x2, 8  -> 1 != ffff -> 참 (다음 조건문으로 바로 감.)
            // rom[5] = 32'b00000000000000000000_00011_0010111; //AUIPC x3 0 -> RF[3] = PC (0x14)
            // rom[6] = 32'b0_000000_00010_00001_100_0100_0_1100011; //BLT x1, x2, 8  -> (signed) 1 < ffff -> 거짓 (다음에 값 나옴)
            // rom[7] = 32'b00000000000000000000_00011_0010111; //AUIPC x3 0 -> RF[3] = PC (0x14)
            // rom[8] = 32'b0_000000_00010_00001_101_0100_0_1100011; //BGE x1, x2, 8  -> (signed) 1 >= ffff -> 참 (다음 조건 문으로 넘어감)
            // rom[9] = 32'b00000000000000000000_00011_0010111; //AUIPC x3 0 -> RF[3] = PC (0x14)
            // rom[10] = 32'b0_000000_00010_00001_110_0100_0_1100011; //BLTU x1, x2, 8 -> (unsigned) 1 < ffff -> 참 (다음 조건문 넘어감)
            // rom[11] = 32'b00000000000000000000_00011_0010111; //AUIPC x3 0 -> RF[3] = PC (0x14)
            // rom[12] = 32'b0_000000_00010_00001_111_0100_0_1100011; //BGEU x1, x2, 8 -> (unsigned) 1 >= ffff -> 거짓 (다음 조건문으로 넘어감)
            // rom[13] = 32'b00000000000000000000_00011_0010111; //AUIPC x3 0 -> RF[3] = PC (0x14)
          
          // U-type test
            // rom[0] = 32'h000010b7; // LUI x1 = 1 << 12
            // rom[1] = 32'h00001117; // AUIPC x2 = PC + (1<<12)
            
            // 0_000 ADD
            // 1_000 SUB
            // 0_001 SLL
            // 0_101 SRL
            // 1_101 SRA
            // 0_010 SLT
            // 0_011 SLTU
            // 0_100 XOR
            // 0_110 OR
            // 0_111 AND


          //main test
          // rom[0]=32'hfe010113;
          // rom[1]=32'h00112e23;
          // rom[2]=32'h00812c23;
          // rom[3]=32'h02010413;
          // rom[4]=32'h00a00793;
          // rom[5]=32'hfef42623;
          // rom[6]=32'h01400793;
          // rom[7]=32'hfef42423;
          // rom[8]=32'hfec42703;
          // rom[9]=32'hfe842783;
          // rom[10]=32'h00f707b3;
          // rom[11]=32'hfef42223;
          // rom[12]=32'hfe442783;
          // rom[13]=32'h00079a63;
          // rom[14]=32'hfec42703;
          // rom[15]=32'hfe842783;
          // rom[16]=32'h40f707b3;
          // rom[17]=32'hfef42223;
          // rom[18]=32'hfec42783;
          // rom[19]=32'hfef42223;
          // rom[20]=32'hfe842583;
          // rom[21]=32'hfec42503;
          // rom[22]=32'h020000ef;
          // rom[23]=32'hfea42423;
          // rom[24]=32'h00000793;
          // rom[25]=32'h00078513;
          // rom[26]=32'h01c12083;
          // rom[27]=32'h01812403;
          // rom[28]=32'h02010113;
          // rom[29]=32'h00008067;
          // rom[30]=32'hfe010113;
          // rom[31]=32'h00812e23;
          // rom[32]=32'h02010413;
          // rom[33]=32'hfea42623;
          // rom[34]=32'hfeb42423;
          // rom[35]=32'hfe842783;
          // rom[36]=32'h4017d793; // rom[36]=32'h0017d793;
          // rom[37]=32'hfef42423;
          // rom[38]=32'hfe842783;
          // rom[39]=32'h00078513;
          // rom[40]=32'h01c12403;
          // rom[41]=32'h02010113;
          // rom[42]=32'h00008067;

        
       

    end

    assign data = rom[addr[31:2]];
endmodule
